Hello! This is an first attempt to creat something
